package PkgUtilities is
  
  type CoreOperation_t is (NoOperation, ForwardPass, BackwardPass);
  
end package PkgUtilities;

package body PkgUtilities is
  
end package body PkgUtilities;
